module vlog_params
  (foo, bar);

  parameter PARAM1 = 1, PARAM2 = 2;

  input wire foo;
  output reg bar;
endmodule;
